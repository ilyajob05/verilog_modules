`timescale 1ns / 1ps

module buttonTest;

	// Inputs
	reg btn1;
	reg btn2;
	reg btn3;
	reg btn4;
	reg clk;
	reg rst;

	// Outputs
	wire led1;
	wire led2;
	wire led3;
	wire led4;

	// Instantiate the Unit Under Test (UUT)
	boardButonLedOnOff uut (
		.btn1(btn1), 
		.btn2(btn2), 
		.btn3(btn3), 
		.btn4(btn4), 
		.led1(led1), 
		.led2(led2), 
		.led3(led3), 
		.led4(led4), 
		.clk(clk), 
		.nrst(rst)
	);

	initial begin
		// Initialize Inputs
		btn1 = 0;
		btn2 = 0;
		btn3 = 0;
		btn4 = 0;
		clk = 0;
		rst = 0;

		// Wait 100 ns for global reset to finish
		#50;
      rst = 1;
		#50;
		// Add stimulus here
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#50;
		btn1 = 1;
		#10;
		btn1 = 0;
		#33;
		btn1 = 1;
		#10;
		btn1 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn1 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#50;
		btn1 = 1;
		#10;
		btn1 = 0;
		#33;
		btn1 = 1;
		#10;
		btn1 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn1 = 0;
		#500;
		
		
		
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#50;
		btn1 = 1;
		#10;
		btn1 = 0;
		#33;
		btn1 = 1;
		#10;
		btn1 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn1 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#10;
		btn1 = 1;
		#10;
		btn1 = 0;
		#50;
		btn1 = 1;
		#10;
		btn1 = 0;
		#33;
		btn1 = 1;
		#10;
		btn1 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn1 = 0;
		#500;
		
		
		
		//кнопка 2 //////////////////////////////
				// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#50;
		btn2 = 1;
		#10;
		btn2 = 0;
		#33;
		btn2 = 1;
		#10;
		btn2 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn2 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#50;
		btn2 = 1;
		#10;
		btn2 = 0;
		#33;
		btn2 = 1;
		#10;
		btn2 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn2 = 0;
		#500;
		
		
		
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#50;
		btn2 = 1;
		#10;
		btn2 = 0;
		#33;
		btn2 = 1;
		#10;
		btn2 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn2 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#10;
		btn2 = 1;
		#10;
		btn2 = 0;
		#50;
		btn2 = 1;
		#10;
		btn2 = 0;
		#33;
		btn2 = 1;
		#10;
		btn2 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn2 = 0;
		#500;
		
		
		//кнопка 3 ///////////////////////////////////////////////////////////////////////////////
				// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#50;
		btn3 = 1;
		#10;
		btn3 = 0;
		#33;
		btn3 = 1;
		#10;
		btn3 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn3 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#50;
		btn3 = 1;
		#10;
		btn3 = 0;
		#33;
		btn3 = 1;
		#10;
		btn3 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn3 = 0;
		#500;
		
		
		
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#50;
		btn3 = 1;
		#10;
		btn3 = 0;
		#33;
		btn3 = 1;
		#10;
		btn3 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn3 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#10;
		btn3 = 1;
		#10;
		btn3 = 0;
		#50;
		btn3 = 1;
		#10;
		btn3 = 0;
		#33;
		btn3 = 1;
		#10;
		btn3 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn3 = 0;
		#500;
		
		
		// кнопка 4 ////////////////////////////////////////////////////////////////////////////////
				// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#50;
		btn4 = 1;
		#10;
		btn4 = 0;
		#33;
		btn4 = 1;
		#10;
		btn4 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn4 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#50;
		btn4 = 1;
		#10;
		btn4 = 0;
		#33;
		btn4 = 1;
		#10;
		btn4 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn4 = 0;
		#500;
		
		
		
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#50;
		btn4 = 1;
		#10;
		btn4 = 0;
		#33;
		btn4 = 1;
		#10;
		btn4 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////
		
		//включение кнопки
		btn4 = 1;
		#500;
		
		// эмуляция дребезга, длительность < 10 ///////////////////////////////////////////
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#10;
		btn4 = 1;
		#10;
		btn4 = 0;
		#50;
		btn4 = 1;
		#10;
		btn4 = 0;
		#33;
		btn4 = 1;
		#10;
		btn4 = 0;
		#77;
		///////////////////////////////////////////////////////////////////////////////////////

		//выключение кнопки
		btn1 = 0;
		#500;
		

	end
      
		
		always #1
			clk <= ~clk;
		
		
endmodule
